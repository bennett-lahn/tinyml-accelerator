// rtl/sys_types.svh
`ifndef SYS_TYPES_SVH
`define SYS_TYPES_SVH
  typedef logic signed [7:0]   int8_t;
  typedef logic signed [15:0] int16_t;
  typedef logic signed [31:0] int32_t;
`endif
